module and_operator(R,A,B);
input [31:0] A;
input [31:0] B;
output [31:0] R;

and (R[0],A[0],B[0]);
and (R[1],A[1],B[1]);
and (R[2],A[2],B[2]);
and (R[3],A[3],B[3]);
and (R[4],A[4],B[4]);
and (R[5],A[5],B[5]);
and (R[6],A[6],B[6]);
and (R[7],A[7],B[7]);
and (R[8],A[8],B[8]);
and (R[9],A[9],B[9]);
and (R[10],A[10],B[10]);
and (R[11],A[11],B[11]);
and (R[12],A[12],B[12]);
and (R[13],A[13],B[13]);
and (R[14],A[14],B[14]);
and (R[15],A[15],B[15]);
and (R[16],A[16],B[16]);
and (R[17],A[17],B[17]);
and (R[18],A[18],B[18]);
and (R[19],A[19],B[19]);
and (R[20],A[20],B[20]);
and (R[21],A[21],B[21]);
and (R[22],A[22],B[22]);
and (R[23],A[23],B[23]);
and (R[24],A[24],B[24]);
and (R[25],A[25],B[25]);
and (R[26],A[26],B[26]);
and (R[27],A[27],B[27]);
and (R[28],A[28],B[28]);
and (R[29],A[29],B[29]);
and (R[30],A[30],B[30]);
and (R[31],A[31],B[31]);

endmodule
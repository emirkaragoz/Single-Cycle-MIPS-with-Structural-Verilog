module nor_operator(R,A,B);
input [31:0] A;
input [31:0] B;
output [31:0] R;

nor (R[0],A[0],B[0]);
nor (R[1],A[1],B[1]);
nor (R[2],A[2],B[2]);
nor (R[3],A[3],B[3]);
nor (R[4],A[4],B[4]);
nor (R[5],A[5],B[5]);
nor (R[6],A[6],B[6]);
nor (R[7],A[7],B[7]);
nor (R[8],A[8],B[8]);
nor (R[9],A[9],B[9]);
nor (R[10],A[10],B[10]);
nor (R[11],A[11],B[11]);
nor (R[12],A[12],B[12]);
nor (R[13],A[13],B[13]);
nor (R[14],A[14],B[14]);
nor (R[15],A[15],B[15]);
nor (R[16],A[16],B[16]);
nor (R[17],A[17],B[17]);
nor (R[18],A[18],B[18]);
nor (R[19],A[19],B[19]);
nor (R[20],A[20],B[20]);
nor (R[21],A[21],B[21]);
nor (R[22],A[22],B[22]);
nor (R[23],A[23],B[23]);
nor (R[24],A[24],B[24]);
nor (R[25],A[25],B[25]);
nor (R[26],A[26],B[26]);
nor (R[27],A[27],B[27]);
nor (R[28],A[28],B[28]);
nor (R[29],A[29],B[29]);
nor (R[30],A[30],B[30]);
nor (R[31],A[31],B[31]);

endmodule